module inversor_8bits (
    input  [7:0] entrada,
    output [7:0] saida
);

    not (saida[0], entrada[0]);
    not (saida[1], entrada[1]);
    not (saida[2], entrada[2]);
    not (saida[3], entrada[3]);
    not (saida[4], entrada[4]);
    not (saida[5], entrada[5]);
    not (saida[6], entrada[6]);
    not (saida[7], entrada[7]);

endmodule